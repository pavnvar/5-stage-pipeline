`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    01:50:22 02/13/2024 
// Design Name: 
// Module Name:    1bit_FS 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module 1bit_FS(
    input A,
    input B,
    input Bin,
    output Out,
    output Bout
    );


endmodule
