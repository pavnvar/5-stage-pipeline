`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    02:23:45 02/13/2024 
// Design Name: 
// Module Name:    fs_64_bit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module fs_64_bit(
    input [63:0] A,
    input [63:0] B,
    input Bin,
    output Bout,
    output [63:0] Diff
    );


endmodule
